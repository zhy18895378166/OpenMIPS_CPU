`include "rtl/include/defines.v"

//时间单位是1ns，精度1ps
`timescale			1ns/1ps

module openmips_min_sopc_tb();

	reg			clock;
	reg			rst;
	
/************************************************************************************************/
/*										第一段：(clk)生成时钟信号									*/
/************************************************************************************************/	
	//每隔10ns，clock翻转一次，所有T=20ns， f= 50MHz
	initial begin
		clock = 1'b0;
		forever #10  clock = ~clock;
	end
	
/************************************************************************************************/
/*										第二段：(rst)复位信号控制									*/
/************************************************************************************************/		
	//最初时刻，复位信号有效，在第195ns，复位信号无效，最小SOPC开始运行
	//在1000ns时，暂停仿真
	initial begin
		rst		= `RstEnable;
		#195 	rst = `RstDisable;
		#1000	$stop;
	end
	
/************************************************************************************************/
/*										第三段：例化最小SOPC									*/
/************************************************************************************************/
	
	//例化指令存储器ROM
	openmips_min_sopc openmips_min_sopc0(
		.clk(clock),
		.rst(rst)
	);
	
endmodule